library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
library ice;
use ice.all;
entity program_memory  is  

port (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(17 DOWNTO 0)
  );
end program_memory;  

architecture Behavioral of program_memory is
component SB_RAM2048x2 is
	generic ( 
       INIT_0 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_1 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_2 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_3 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_4 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_5 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_6 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_7 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_8 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_9 : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_A : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_B : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_C : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_D : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_E : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
       INIT_F : bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
       ) ;
      port( 
          RDATA : out std_logic_vector( 1  downto 0) ;
          RCLK  : in  std_logic ;
          RCLKE : in  std_logic := 'H';
          RE    : in  std_logic := 'L';
          RADDR : in  std_logic_vector( 10  downto 0) ;
          WCLK  : in  std_logic ;
          WCLKE : in  std_logic := 'H';
          WE    : in  std_logic := 'L';
          WADDR : in  std_logic_vector( 10  downto 0) ;
          WDATA : in  std_logic_vector( 1  downto 0)
         );
end component;
signal WE : std_logic;
begin 
WE <= wea(0);
Ram2048x2_inst0 : SB_RAM2048x2
generic map (
INIT_0 => X"0020303259393935E44E4E493B46011C140140EBF2DDB402EC845046384100511",
INIT_1 => X"13417414100100442221220055D1D891E0005591E8D1D052200444098A072A001",
INIT_2 => X"1430074685C4074685C44194CBC2F48C1027C000019230939384E4E4E4E848393",
INIT_3 => X"3939320008C048393939325E429393219394E4E80000C248F4E429393540E5300",
INIT_4 => X"00C4119411650C01C1000170000140E49300C32DC4F384135300000AAA2000094",
INIT_5 => X"4FF3A00084C6C60E429835E01939B49315E4224E4E6A500B50240409000000204",
INIT_6 => X"46444458C42A39F4210117644409C0426E4E49342E939BAAA644444440906939B",
INIT_7 => X"BAAA4444454265E4AAAA8888090A5E4AAAAA8888948AAA0000E429C8AAA0000E4",
INIT_8 => X"493010110008180490C1818D8829CF3A080022088001200800320802000520240",
INIT_9 => X"000848054A90F9E493101728394414D914E4A000200802008120000C0C6C60000",
INIT_A => X"083944E4E4930E497460005935E4E4E4930200000094E4E49335E000035E09394",
INIT_B => X"4E420004E4A35E100835E51200411839C3127400142033218C04E4E01FF800208",
INIT_C => X"88002204800020C80080004100000000000000000000000000000000000000000",
INIT_D => X"00000000000000000000000000000000000000000000000000000000000000000",
INIT_E => X"00000000000000000000000000000000000000000000000000000000000000000",
INIT_F => X"00000000000000000000000000000000000000000000000000000000000000000"
)
port map (
RDATA => douta(1 downto 0),
RADDR => addra(10 downto 0),
RCLK => clka,
RCLKE => ena,
RE => '1',
WADDR => addra(10 downto 0),
WCLK=> clka,
WCLKE => ena,
WDATA => dina(1 downto 0),
WE => WE
);
Ram2048x2_inst1 : SB_RAM2048x2
generic map (
INIT_0 => X"55000A0460004592050055A044146090649545000441454100500854155242201",
INIT_1 => X"11A0000000980028888888A055424640488055404642480110600400010001014",
INIT_2 => X"40010505050544444444440001694040121000000019000451400550055402451",
INIT_3 => X"1045112004600045104519205104519A045005548008058012051045125054100",
INIT_4 => X"004849504002042849AAA04AAA22145A040940011448445051000005551000014",
INIT_5 => X"41115000444510005104920100451A04920555005500010140181100000000102",
INIT_6 => X"25666A000010451510220856666104811055A0001104555555666201014010455",
INIT_7 => X"5555101010A11205555510008605205555500000044555000005104455500005A",
INIT_8 => X"A0401119AAA40440001440405454455150190842029284202918442100041015A",
INIT_9 => X"AAA604015101015A0050540045002021000550001004610040100002045100000",
INIT_A => X"004500055A0405A0415AAA049200055A044100000040055A04920100092010450",
INIT_B => X"005100000559209AA692000100841400010100440998001042000550055551442",
INIT_C => X"2029084A029084602140000100000000000000000000000000000000000000000",
INIT_D => X"00000000000000000000000000000000000000000000000000000000000000000",
INIT_E => X"00000000000000000000000000000000000000000000000000000000000000000",
INIT_F => X"00000000000000000000000000000000000000000000000000000000000000000"
)
port map (
RDATA => douta(3 downto 2),
RADDR => addra(10 downto 0),
RCLK => clka,
RCLKE => ena,
RE => '1',
WADDR => addra(10 downto 0),
WCLK=> clka,
WCLKE => ena,
WDATA => dina(3 downto 2),
WE => WE
);
Ram2048x2_inst2 : SB_RAM2048x2
generic map (
INIT_0 => X"0000101ABF30000000555555521387045C17D901304AAAEA05CAAA8EA8A203103",
INIT_1 => X"31000C0601CC4034DDFCDDC4008E638F7F0500CC430C4F023040050013C043040",
INIT_2 => X"000049494949494949490AFDD7C2E2E92056900081A6A05555800005555800004",
INIT_3 => X"4555120404401000455512000455512000055558001003046000455515AE04593",
INIT_4 => X"390696AF4031833E40000030008B28AAAA66421298424852615E424AAAB000028",
INIT_5 => X"844C20000855551559A8AAA2000080000000880000EFB20400949128000000201",
INIT_6 => X"130004D45001004592022230008ECD002008AA20BF0000AAA2000CCDC1CA70000",
INIT_7 => X"0AAACDDEDC0BB0000AAADCCC0CAF0000AAAFDCECC49AAE2000559A49AAE2000AA",
INIT_8 => X"AAA89800000B0B2DF1C0B0BC832C300A0980421490052389806219700008E1E00",
INIT_9 => X"00083838AAF19DAAAAA1A63755A6549D100000000000400000000029165551000",
INIT_A => X"0455A55555550AAAE120000AAAA55555558000000005555555000C49300000005",
INIT_B => X"555D4930008AAA0008AAA0100049AB0FDBB7202150316A3189245551800824210",
INIT_C => X"09005234980621890410000200000000000000000000000000000000000000000",
INIT_D => X"00000000000000000000000000000000000000000000000000000000000000000",
INIT_E => X"00000000000000000000000000000000000000000000000000000000000000000",
INIT_F => X"00000000000000000000000000000000000000000000000000000000000000000"
)
port map (
RDATA => douta(5 downto 4),
RADDR => addra(10 downto 0),
RCLK => clka,
RCLKE => ena,
RE => '1',
WADDR => addra(10 downto 0),
WCLK=> clka,
WCLKE => ena,
WDATA => dina(5 downto 4),
WE => WE
);
Ram2048x2_inst3 : SB_RAM2048x2
generic map (
INIT_0 => X"00804040000000000000000004400080008000000400000400400000400004004",
INIT_1 => X"40008000080000400000000000000400000000040404000400080000440000000",
INIT_2 => X"04000000000000000000040004000000004000000004080000000000000000000",
INIT_3 => X"00000400000008000000040000000040000000000008008000000000000000000",
INIT_4 => X"00000000000000000000000000000000000000000844000400800000004000000",
INIT_5 => X"00000000080000000000000000000000000000000000000000004440080000400",
INIT_6 => X"04000008000000000000004000008000000000000000000004000048880000000",
INIT_7 => X"00008080800040000000040800040000000000000000000000000000000000000",
INIT_8 => X"00000000000000000080000080004000000404000040400004040040000000080",
INIT_9 => X"00000000000000000000040000040000400040000000000000000040040000000",
INIT_A => X"00000000000000000000000000000000000000000000000000000000000000000",
INIT_B => X"00000000004000000000000000000000040000004044000400000000000000400",
INIT_C => X"00040400004040000000000000000000000000000000000000000000000000000",
INIT_D => X"00000000000000000000000000000000000000000000000000000000000000000",
INIT_E => X"00000000000000000000000000000000000000000000000000000000000000000",
INIT_F => X"00000000000000000000000000000000000000000000000000000000000000000"
)
port map (
RDATA => douta(7 downto 6),
RADDR => addra(10 downto 0),
RCLK => clka,
RCLKE => ena,
RE => '1',
WADDR => addra(10 downto 0),
WCLK=> clka,
WCLKE => ena,
WDATA => dina(7 downto 6),
WE => WE
);
Ram2048x2_inst4 : SB_RAM2048x2
generic map (
INIT_0 => X"00818100000000000000000009C010460140100114555555555555555555A4990",
INIT_1 => X"0B23400EE01181421111111C55144C3CC10D55144C3CC11004172089DA876A455",
INIT_2 => X"5A516363636363636363CE956D7F55665995611199566100048B1B1B1B18B6C6C",
INIT_3 => X"C6C60644554CB6C6C6C60E6C6C6C60EA1B1B1B18115D57B566C6C6C601B4A86E4",
INIT_4 => X"4E86CA60840A394296C614A1B50A296C6900802CB0B280E282939F29393939380",
INIT_5 => X"08801111D75E4E1B1B181B50C6C606C6D6C6B06C6D66A34890A8262809393F238",
INIT_6 => X"8FEEEE2CC8A6C64C60F338FEEEE2CC8A6C64C60BBF6C681B174440030FEAF6C68",
INIT_7 => X"81B1303030BBF6C691B53000CEAF6C691B530000084E4E4E4EB1B18493949396C",
INIT_8 => X"C61C088B1B1444036A004440852D0081111644811164481116448544E4E1141C6",
INIT_9 => X"6C64050B7298016C649994881B1566211C6CA393E4E00E4E04444406A93931C61",
INIT_A => X"1B1B1C61B1B166C68191B1991B1C61B1B154E4E4935C61B1B1C6139396C60B5C6",
INIT_B => X"6C609396C681B16C681B161E4E4C2119559955669510999989500001100664481",
INIT_C => X"11164481116448111619397200000000000000000000000000000000000000000",
INIT_D => X"00000000000000000000000000000000000000000000000000000000000000000",
INIT_E => X"00000000000000000000000000000000000000000000000000000000000000000",
INIT_F => X"00000000000000000000000000000000000000000000000000000000000000000"
)
port map (
RDATA => douta(9 downto 8),
RADDR => addra(10 downto 0),
RCLK => clka,
RCLKE => ena,
RE => '1',
WADDR => addra(10 downto 0),
WCLK=> clka,
WCLKE => ena,
WDATA => dina(9 downto 8),
WE => WE
);
Ram2048x2_inst5 : SB_RAM2048x2
generic map (
INIT_0 => X"00000000000000000000000000000040080080044000000000000000000000000",
INIT_1 => X"00440000004404004444444000400040040000400040040800800800000000000",
INIT_2 => X"00040404040404040404000000000000000000008004000000000000000000400",
INIT_3 => X"00400008088000400040000400040000000000000000040840400040000000000",
INIT_4 => X"00000040400000000040000000000004080800000000000000000000004000080",
INIT_5 => X"04400000048000800000000800400040004000040000400880000008000040000",
INIT_6 => X"00000040000040040000000000040000040040000404000000000800000040400",
INIT_7 => X"00000000000040400000000000040400000000000000000000000000000000004",
INIT_8 => X"40004000000000000000000040000080000044800004480000448000000000000",
INIT_9 => X"04000080000400040000004000000000400400000000000000000000000000400",
INIT_A => X"00000400000000400400000000040000000000000004000000400400004000000",
INIT_B => X"04000000400000040000004000800000004000004000000000000000000004480",
INIT_C => X"00004480000448000080000400000000000000000000000000000000000000000",
INIT_D => X"00000000000000000000000000000000000000000000000000000000000000000",
INIT_E => X"00000000000000000000000000000000000000000000000000000000000000000",
INIT_F => X"00000000000000000000000000000000000000000000000000000000000000000"
)
port map (
RDATA => douta(11 downto 10),
RADDR => addra(10 downto 0),
RCLK => clka,
RCLKE => ena,
RE => '1',
WADDR => addra(10 downto 0),
WCLK=> clka,
WCLKE => ena,
WDATA => dina(11 downto 10),
WE => WE
);
Ram2048x2_inst6 : SB_RAM2048x2
generic map (
INIT_0 => X"AA45454AAAAAAAAAAAAAAAAAA5020205014010888655555555555555555512596",
INIT_1 => X"658569659611144B1111111100466C46605100466C46605461157750435003501",
INIT_2 => X"1564525252525252525210A88A82A888222A800002A9A7AAAA5AAAAAAAA5A9AAA",
INIT_3 => X"AAAA69E3A89988AAAAAA69AAAAAAA696AAAAAAA5AF8A8B98B9AAAAAA6AA793C55",
INIT_4 => X"5578AAAA8D2639851000092000066AAAAACA8262890A890620AAA2EFFF7FFF7A9",
INIT_5 => X"90082000C88AAA6AAAA9AAA6BAAAAAAAAAAAAAAAAAAA2C5491A822695CFF7266A",
INIT_6 => X"A30008A8993AAAAAA6266A30008A8993AAAAAA6A3AAAA2AAA200089A9AE3AAAA2",
INIT_7 => X"2AAAA9A9A9A3AAAA2AAAA9999E3AAAA2AAAA999991FFFFDFFFAAAA1FFFFDFFFAA",
INIT_8 => X"AAA12660000ADA88A2A8ADA9A2AD00088810260881026088102600200009A8A20",
INIT_9 => X"00086B6008A228AAA2A8A02AAAA82A284AAA2000000C8000CD00003AE8AAA6555",
INIT_A => X"59AAAAAAAAAA5AAA2220005AAAAAAAAAAA800000009AAAAAAAAAA2AAAAAAAAAAA",
INIT_B => X"AAAAAAAAAAAAAA0008AAA560008A266A8222A8882A9A22265AE9AAA6100022608",
INIT_C => X"88102608810260881000004600000000000000000000000000000000000000000",
INIT_D => X"00000000000000000000000000000000000000000000000000000000000000000",
INIT_E => X"00000000000000000000000000000000000000000000000000000000000000000",
INIT_F => X"00000000000000000000000000000000000000000000000000000000000000000"
)
port map (
RDATA => douta(13 downto 12),
RADDR => addra(10 downto 0),
RCLK => clka,
RCLKE => ena,
RE => '1',
WADDR => addra(10 downto 0),
WCLK=> clka,
WCLKE => ena,
WDATA => dina(13 downto 12),
WE => WE
);
Ram2048x2_inst7 : SB_RAM2048x2
generic map (
INIT_0 => X"00000000000000000000000000040000000000040000000000000000000000080",
INIT_1 => X"00080400800004000000000400400040004000400040000404040000000000400",
INIT_2 => X"00400000000000000000400400400400000400000040000000400000000404000",
INIT_3 => X"00000000040044000000000000000000000000040004004004000000000004000",
INIT_4 => X"00000004000400000000080000000000044440040000400040000000004000040",
INIT_5 => X"00000000440000000004000040000000000000000040404400440000000000404",
INIT_6 => X"40000040000400000004040000040000400000000000000000000400000000000",
INIT_7 => X"00000000000000000000404040000000000004040400000000000040000000000",
INIT_8 => X"00000000000000440000000000400044400000040000004000000000000008000",
INIT_9 => X"00040000040040000008000400000040000000000004400040000000400000000",
INIT_A => X"00000000000000000000000000000000004000000000000000000000000040000",
INIT_B => X"00000000004000000000000000400000400044000400000440400000000000004",
INIT_C => X"40000004000000400000000000000000000000000000000000000000000000000",
INIT_D => X"00000000000000000000000000000000000000000000000000000000000000000",
INIT_E => X"00000000000000000000000000000000000000000000000000000000000000000",
INIT_F => X"00000000000000000000000000000000000000000000000000000000000000000"
)
port map (
RDATA => douta(15 downto 14),
RADDR => addra(10 downto 0),
RCLK => clka,
RCLKE => ena,
RE => '1',
WADDR => addra(10 downto 0),
WCLK=> clka,
WCLKE => ena,
WDATA => dina(15 downto 14),
WE => WE
);
Ram2048x2_inst8 : SB_RAM2048x2
generic map (
INIT_0 => X"AA20202AAAAAAAAAAAAAAAAAA02BAAA0A82A8AEDDAAAAAAAAAAAAAAAAAAA0B05B",
INIT_1 => X"B0CD2AA05B88AD698888888255D662D6682055D662D6685CA2965D2A082A28228",
INIT_2 => X"843A0808080808080808AA0CC2C0BCCC233BC55513B000AAAA20000AAAA200008",
INIT_3 => X"8AAAA0000C8000008AAAA00008AAAA00000AAAA20000C80C80008AAAA005FB655",
INIT_4 => X"55F200A2C5075D538555557555136DAAA202C03AA8A2C8A2A65551300045551A8",
INIT_5 => X"8AA24555108AAAA000020008300000008AAA0AAAAA28AE2D92BC2338055590322",
INIT_6 => X"2455592C8002008AAA0322455592C8002008AAA00C000000075551828204D0000",
INIT_7 => X"000038282800C00000003828204D0000000382828A00005555AAAAA00005555AA",
INIT_8 => X"AAA2332555505A8C003C05A820C0459CD916768D916768D916768135555D05A65",
INIT_9 => X"555149AAAD03BA000805AA23000249AAA00045555551C5551555550008AAAA000",
INIT_A => X"00000AAAAAAA00004375555AAAA0000000D5555555DAAAAAAA0004555AAA20000",
INIT_B => X"0004555AAA20005559AAA1A555104590C233BCCC2B0823332008AAAA05527768D",
INIT_C => X"D916768D916768D91645555B00000000000000000000000000000000000000000",
INIT_D => X"00000000000000000000000000000000000000000000000000000000000000000",
INIT_E => X"00000000000000000000000000000000000000000000000000000000000000000",
INIT_F => X"00000000000000000000000000000000000000000000000000000000000000000"
)
port map (
RDATA => douta(17 downto 16),
RADDR => addra(10 downto 0),
RCLK => clka,
RCLKE => ena,
RE => '1',
WADDR => addra(10 downto 0),
WCLK=> clka,
WCLKE => ena,
WDATA => dina(17 downto 16),
WE => WE
);
end Behavioral;

